module data(
    input       [2:0]   pulse,
    input       [5:0]   seq,
    output              e,
    output  reg         rs,
                        rw,
    output  reg [3:0]   note,
    output  reg [7:0]   disp_c_n,
                        disp_s,
                        db,
    output  reg [63:0]  col_r_data,
                        col_g_data
);
///////////////////////////////////////////////
    always @(*)
        case (seq)
            6'd2: begin
                col_r_data  =
                {
                    8'b0000_0000,
                    8'b0001_0000,
                    8'b0010_1000,
                    8'b0011_1000,
                    8'b0000_1000,
                    8'b0011_0000,
                    8'b0000_0000,
                    8'b0000_0000
                };
                col_g_data  =
                {
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0100,
                    8'b0001_0100,
                    8'b0000_0100,
                    8'b0001_1000,
                    8'b0000_0000
                };
            end
            6'd3: begin
                col_r_data  =
                {
                    8'b0000_0000,
                    8'b0001_0000,
                    8'b0010_1000,
                    8'b0011_1000,
                    8'b0010_1000,
                    8'b0001_0000,
                    8'b0000_0000,
                    8'b0000_0000
                };
                col_g_data  =
                {
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0100,
                    8'b0001_0100,
                    8'b0000_0100,
                    8'b0000_1000,
                    8'b0000_0000
                };
            end
            6'd4: begin
                col_r_data  =
                {
                    8'b0000_0000,
                    8'b0011_1000,
                    8'b0010_1000,
                    8'b0000_1000,
                    8'b0001_0000,
                    8'b0001_0000,
                    8'b0000_0000,
                    8'b0000_0000
                };
                col_g_data  =
                {
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0001_0100,
                    8'b0001_0100,
                    8'b0000_0100,
                    8'b0000_1000,
                    8'b0000_1000,
                    8'b0000_0000
                };
            end
            6'd5: begin
                col_r_data  =
                {
                    8'b0000_0000,
                    8'b0001_1000,
                    8'b0010_0000,
                    8'b0011_1000,
                    8'b0010_1000,
                    8'b0001_0000,
                    8'b0000_0000,
                    8'b0000_0000
                };
                col_g_data  =
                {
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_1100,
                    8'b0000_0000,
                    8'b0001_0100,
                    8'b0000_0100,
                    8'b0000_1000,
                    8'b0000_0000
                };
            end
            6'd6: begin
                col_r_data  =
                {
                    8'b0000_0000,
                    8'b0011_1000,
                    8'b0010_0000,
                    8'b0001_0000,
                    8'b0000_1000,
                    8'b0011_1000,
                    8'b0000_0000,
                    8'b0000_0000
                };
                col_g_data  =
                {
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0001_1100,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0100,
                    8'b0001_1100,
                    8'b0000_0000
                };
            end
            6'd7: begin
                col_r_data  =
                {
                    8'b0000_0000,
                    8'b0001_1000,
                    8'b0010_1000,
                    8'b0010_1000,
                    8'b0011_1100,
                    8'b0000_1000,
                    8'b0000_0000,
                    8'b0000_0000
                };
                col_g_data  =
                {
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0100,
                    8'b0000_0100,
                    8'b0000_0000,
                    8'b0001_0110,
                    8'b0000_0100,
                    8'b0000_0000
                };
            end
            6'd8: begin
                col_r_data  =
                {
                    8'b0000_0000,
                    8'b0011_0000,
                    8'b0000_1000,
                    8'b0001_0000,
                    8'b0000_1000,
                    8'b0011_0000,
                    8'b0000_0000,
                    8'b0000_0000
                };
                col_g_data  =
                {
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0001_0000,
                    8'b0000_0100,
                    8'b0000_0000,
                    8'b0000_0100,
                    8'b0001_1000,
                    8'b0000_0000
                };
            end
            6'd9: begin
                col_r_data  =
                {
                    8'b0000_0000,
                    8'b0001_0000,
                    8'b0010_1000,
                    8'b0000_1000,
                    8'b0001_0000,
                    8'b0011_1000,
                    8'b0000_0000,
                    8'b0000_0000
                };
                col_g_data  =
                {
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0001_0100,
                    8'b0000_0100,
                    8'b0000_0000,
                    8'b0001_1100,
                    8'b0000_0000
                };
            end
            6'd10: begin
                col_r_data  =
                {
                    8'b0000_0000,
                    8'b0001_0000,
                    8'b0011_0000,
                    8'b0001_0000,
                    8'b0001_0000,
                    8'b0011_1000,
                    8'b0000_0000,
                    8'b0000_0000
                };
                col_g_data  =
                {
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_1000,
                    8'b0000_1000,
                    8'b0000_1000,
                    8'b0000_0000,
                    8'b0001_1100,
                    8'b0000_0000
                };
            end
            6'd11: begin
                col_r_data  =
                {
                    8'b0000_0000,
                    8'b0001_0000,
                    8'b0010_1000,
                    8'b0010_1000,
                    8'b0010_1000,
                    8'b0001_0000,
                    8'b0000_0000,
                    8'b0000_0000
                };
                col_g_data  =
                {
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0001_0100,
                    8'b0001_0100,
                    8'b0000_0100,
                    8'b0000_1000,
                    8'b0000_0000
                };
            end
            6'd12:
                case (pulse[2:1])
                    2'd0: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd1: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd2: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0100_0010,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0100_0010,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd3: begin
                        col_r_data  =
                        {
                            8'b1000_0001,
                            8'b0100_0010,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0100_0010,
                            8'b1000_0001
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                endcase
            6'd13:
                case (pulse[2:1])
                    2'd0: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd1: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd2: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0100_0010,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0100_0010,
                            8'b0000_0000
                        };
                    end
                    2'd3: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b1000_0001,
                            8'b0100_0010,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0100_0010,
                            8'b1000_0001
                        };
                    end
                endcase
            6'd14:
                case (pulse[2:1])
                    2'd0: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd1: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd2: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0100_0010,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0100_0010,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0100_0010,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0100_0010,
                            8'b0000_0000
                        };
                    end
                    2'd3: begin
                        col_r_data  =
                        {
                            8'b1000_0001,
                            8'b0100_0010,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0100_0010,
                            8'b1000_0001
                        };
                        col_g_data  =
                        {
                            8'b1000_0001,
                            8'b0100_0010,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0100_0010,
                            8'b1000_0001
                        };
                    end
                endcase
            6'd15:
                case (pulse[2:1])
                    2'd0: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd1: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd2: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0011_1100,
                            8'b0100_0010,
                            8'b0100_0010,
                            8'b0100_0010,
                            8'b0100_0010,
                            8'b0011_1100,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd3: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0111_1110,
                            8'b1000_0001,
                            8'b1000_0001,
                            8'b1000_0001,
                            8'b1000_0001,
                            8'b1000_0001,
                            8'b1000_0001,
                            8'b0111_1110
                        };
                    end
                endcase
            6'd16:
                case (pulse[2:1])
                    2'd0: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd1: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd2: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0011_1100,
                            8'b0100_0010,
                            8'b0100_0010,
                            8'b0100_0010,
                            8'b0100_0010,
                            8'b0011_1100,
                            8'b0000_0000
                        };
                    end
                    2'd3: begin
                        col_r_data  =
                        {
                            8'b0111_1110,
                            8'b1000_0001,
                            8'b1000_0001,
                            8'b1000_0001,
                            8'b1000_0001,
                            8'b1000_0001,
                            8'b1000_0001,
                            8'b0111_1110
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                endcase
            6'd17:
                case (pulse[2:1])
                    2'd0: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd1: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0010_0100,
                            8'b0010_0100,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd2: begin
                        col_r_data  =
                        {
                            8'b0000_0000,
                            8'b0011_1100,
                            8'b0100_0010,
                            8'b0101_1010,
                            8'b0101_1010,
                            8'b0100_0010,
                            8'b0011_1100,
                            8'b0000_0000
                        };
                        col_g_data  =
                        {
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0001_1000,
                            8'b0001_1000,
                            8'b0000_0000,
                            8'b0000_0000,
                            8'b0000_0000
                        };
                    end
                    2'd3: begin
                        col_r_data  =
                        {
                            8'b0110_1100,
                            8'b0000_0001,
                            8'b1001_1001,
                            8'b1010_0100,
                            8'b0010_0101,
                            8'b1001_1001,
                            8'b1000_0000,
                            8'b0011_0110
                        };
                        col_g_data  =
                        {
                            8'b0011_0110,
                            8'b1000_0000,
                            8'b1000_0001,
                            8'b0000_0001,
                            8'b1000_0000,
                            8'b1000_0001,
                            8'b0000_0001,
                            8'b0110_1100
                        };
                    end
                endcase
            6'd0:
                if (pulse[2] == 1'b0) begin
                    col_r_data  =   {64{1'b0}};
                    col_g_data  =   {64{1'b1}};
                end else begin
                    col_r_data  =   {64{1'b1}};
                    col_g_data  =   {64{1'b0}};
                end
            6'd1:
                if (pulse[2] == 1'b0) begin
                    col_r_data  =   {64{1'b1}};
                    col_g_data  =   {64{1'b1}};
                end else begin
                    col_r_data  =   {64{1'b0}};
                    col_g_data  =   {64{1'b0}};
                end
            default: begin
                col_r_data  =
                {
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000
                };
                col_g_data  =
                {
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000,
                    8'b0000_0000
                };
            end
        endcase
///////////////////////////////////////////////
    parameter off   = 8'b1111_1111;
    parameter on    = 8'b0000_0000;
    parameter on_7  = 8'b0111_1111;

    parameter s_    = 8'b0000_0000;
    parameter s0    = 8'b0011_1111;
    parameter s1    = 8'b0000_0110;
    parameter s2    = 8'b0101_1011;
    parameter s3    = 8'b0100_1111;
    parameter s4    = 8'b0110_0110;
    parameter s5    = 8'b0110_1101;
    parameter s6    = 8'b0111_1101;
    parameter s7    = 8'b0000_0111;
    parameter s8    = 8'b0111_1111;
    parameter s9    = 8'b0110_1111;

    always @(*)
        case (seq)
            6'd2: begin
                    disp_c_n    =   on_7;
                    disp_s      =   s9;
            end
            6'd3: begin
                    disp_c_n    =   on_7;
                    disp_s      =   s8;
            end
            6'd4: begin
                    disp_c_n    =   on_7;
                    disp_s      =   s7;
            end
            6'd5: begin
                    disp_c_n    =   on_7;
                    disp_s      =   s6;
            end
            6'd6: begin
                    disp_c_n    =   on_7;
                    disp_s      =   s5;
            end
            6'd7: begin
                    disp_c_n    =   on_7;
                    disp_s      =   s4;
            end
            6'd8: begin
                    disp_c_n    =   on_7;
                    disp_s      =   s3;
            end
            6'd9: begin
                    disp_c_n    =   on_7;
                    disp_s      =   s2;
            end
            6'd10: begin
                    disp_c_n    =   on_7;
                    disp_s      =   s1;
            end
            6'd11: begin
                    disp_c_n    =   on_7;
                    disp_s      =   s0;
            end
            6'd0:
                if (pulse[1] == 1'b0) begin
                    disp_c_n    =   on;
                    disp_s      =   s8;
                end else begin
                    disp_c_n    =   off;
                    disp_s      =   s_;
                end
            6'd1:
                if (pulse[2:1] == 2'd0) begin
                    disp_c_n    =   on;
                    disp_s      =   s8;
                end else begin
                    disp_c_n    =   off;
                    disp_s      =   s_;
                end
            default: begin
                    disp_c_n    =   off;
                    disp_s      =   s_;
            end
        endcase
///////////////////////////////////////////////
    parameter g  = 4'b0101;
    parameter b  = 4'b0111;
    parameter re = 4'b1000;
    parameter c1 = 4'b1001;
    parameter d1 = 4'b1010;
    parameter e1 = 4'b1011;
    parameter f1 = 4'b1100;
    parameter g1 = 4'b1101;
    parameter a1 = 4'b1110;
    parameter b1 = 4'b1111;
    always @(*)
        case (seq)
            6'd2:
                if (pulse[2:1] == 2'd2)
                            note    =   e1;
                else
                            note    =   d1;
            6'd3:           note    =   c1;
            6'd4:
                if (pulse[2:1] == 2'd2)
                            note    =   e1;
                else
                            note    =   d1;
            6'd5:
                if (pulse[2:0] == 3'd7)
                            note    =   re;
                else
                            note    =   g;
            ////////
            6'd6:
                if (pulse[2] == 1'b0)
                            note    =   g;
                else if (pulse[2:0] == 3'd7)
                            note    =   re;
                else
                            note    =   g1;
            6'd7:
                case (pulse[2:1])
                    2'd0:   note    =   g1;
                    2'd1:   note    =   d1;
                    2'd2:   note    =   f1;
                    2'd3:   note    =   e1;
                endcase
            6'd8:           note    =   d1;
            6'd9:           note    =   d1;
            ////////////////
            6'd10:
                case (pulse[2:1])
                    2'd0:   note    =   b;
                    2'd1:
                        if (pulse[0] == 1'b0)
                            note    =   b;
                        else
                            note    =   c1;
                    2'd2:   note    =   d1;
                    2'd3:   note    =   e1;
                endcase
            6'd11:          note    =   c1;
            6'd12:
                case (pulse[2:1])
                    2'd0:   note    =   b;
                    2'd1:   note    =   c1;
                    2'd2:   note    =   d1;
                    2'd3:   note    =   e1;
                endcase
            6'd13:
                if (pulse[2:0] == 3'd7)
                            note    =   re;
                else
                            note    =   g;
            ////////
            6'd14:
                if (pulse[2] == 1'b0)
                            note    =   g;
                else
                            note    =   f1;
            6'd15:
                case (pulse[2:1])
                    2'd0:   note    =   e1;
                    2'd1:   note    =   f1;
                    2'd2:   note    =   e1;
                    2'd3:   note    =   d1;
                endcase
            6'd16:          note    =   c1;
            6'd17:          note    =   c1;
            ///////////////////////////////
            6'd18:
                if (pulse[2:1] == 2'd2)
                            note    =   a1;
                else
                            note    =   g1;
            6'd19:
                if (pulse[2] == 1'b0)
                            note    =   f1;
                else
                            note    =   c1;
            6'd20:
                case (pulse[2:1])
                    2'd0:   note    =   e1;
                    2'd1:   note    =   f1;
                    2'd2:   note    =   g1;
                    2'd3:   note    =   a1;
                endcase
            6'd21:          note    =   g1;
            ////////
            6'd22:
                if (pulse[2] == 1'b0)
                            note    =   d1;
                else
                            note    =   a1;
            6'd23:
                case (pulse[2:1])
                    2'd0:   note    =   g1;
                    2'd1:   note    =   a1;
                    2'd2:   note    =   f1;
                    2'd3:   note    =   a1;
                endcase
            6'd24:          note    =   g1;
            6'd25:          note    =   g1;
            ////////////////
            6'd26:
                case (pulse[2:1])
                    2'd0:   note    =   e1;
                    2'd1:   note    =   f1;
                    2'd2:   note    =   e1;
                    2'd3:   note    =   d1;
                endcase
            6'd27:          note    =   g;
            6'd28:
                case (pulse[2:1])
                    2'd0:   note    =   e1;
                    2'd1:   note    =   f1;
                    2'd2:   note    =   e1;
                    2'd3:   note    =   d1;
                endcase
            6'd29:          note    =   c1;
            ////////
            6'd30:
                if (pulse[2] == 1'b0)
                            note    =   g;
                else
                            note    =   f1;
            6'd31:
                case (pulse[2:1])
                    2'd0:   note    =   e1;
                    2'd1:   note    =   f1;
                    2'd2:   note    =   e1;
                    2'd3:   note    =   d1;
                endcase
            6'd32:          note    =   c1;
            6'd33:          note    =   re;
            //
            default:        note    =   re;
        endcase
///////////////////////////////////////////////
    // 根据工作状态分配下降沿（写指令使能信号）
    assign e = (seq < 6'd34) ? ((seq < 6'd2) ? ~pulse[0] : ~pulse[2]) : 1'b0;
    parameter idle              = 10'b00_0000_0000; // 空闲，无指令
    parameter function_set      = 10'b00_0011_1000; // Function set
    parameter display_on        = 10'b00_0000_1100; // Display on
    parameter display_clear     = 10'b00_0000_0001; // Display clear
    parameter entry_mode_set    = 10'b00_0000_0110; // Entry mode set
    parameter enter             = 10'b00_1100_0000; // 跳转至40H地址，即第二行
    parameter put_char          = 2'b10;            // 写入数据指令前缀

    wire    [7:0]   char_1  [2:16], // 定义第一行字符地址数据，最多15个字符
                    char_2  [18:32];// 定义第二行字符地址数据，最多15个字符
    assign {
        char_1[2],
        char_1[3],
        char_1[4],
        char_1[5],
        char_1[6],
        char_1[7],
        char_1[8],
        char_1[9],
        char_1[10],
        char_1[11],
        char_1[12],
        char_1[13],
        char_1[14],
        char_1[15],
        char_1[16]
    } = "Happy new year!";          // 装箱第一行字符地址数据
    assign {
        char_2[18],
        char_2[19],
        char_2[20],
        char_2[21],
        char_2[22],
        char_2[23],
        char_2[24],
        char_2[25],
        char_2[26],
        char_2[27],
        char_2[28],
        char_2[29],
        char_2[30],
        char_2[31],
        char_2[32]
    } = "it's near 2020!";          // 装箱第二行字符地址数据

    always @(*)
        if (seq == 6'd0)
                        {rs, rw, db} = function_set;    // 根据datasheet，此处应发送function set指令四次
        else if (seq == 6'd1)
            case (pulse[2:1])
                2'd0:   {rs, rw, db} = display_on;      // 发送display on指令，打开显示
                2'd1:   {rs, rw, db} = {put_char, "*"}; // 向DDRAM写入一个星号对应的地址作为自检测试
                2'd2:   {rs, rw, db} = display_clear;   // 发送display clear指令，清除屏幕，清零地址计数器
                2'd3:   {rs, rw, db} = entry_mode_set;  // 发送entry mode set指令
            endcase                                     // 设置模式为: 地址计数器自动+1, 无光标
        else if (seq >= 6'd2 && seq <= 6'd16)           // 第一行，写入对应地址（与ASCII码一致）
                        {rs, rw, db} = {put_char, char_1[seq]};
        else if (seq == 6'd17)                          // 跳转至第二行开始
                        {rs, rw, db} = enter;
        else if (seq >= 6'd18 && seq <= 6'd32)          // 第二行，写入对应地址（与ASCII码一致）
                        {rs, rw, db} = {put_char, char_2[seq]};
        else if (seq == 6'd33)
                        {rs, rw, db} = display_clear;   // 到达末尾，音乐结束后半秒后清零
        else            {rs, rw, db} = idle;            // 其余情况为空闲

endmodule // data
